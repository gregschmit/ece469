module aludec(input logic [5:0] funct,
              input logic [1:0] aluop,
              output logic [2:0] alucontrol);

 // ADD CODE HERE
 // Complete the design for the ALU Decoder.
 // Your design goes here. Remember that this is a combinational
 // module.
 // Remember that you may also reuse any code from previous labs.
endmodule

